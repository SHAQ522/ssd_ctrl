module ChannelContant(
						output [7 : 0] ch
						);
						
	parameter [7 : 0] ch_p = 8'd0;
	
endmodule 
module clk_df(clk,clk_out);

input clk;
output clk_out;

assign   clk_out = clk;                   


endmodule
